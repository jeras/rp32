////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////

module r5p_tb #(
  // RISC-V ISA
  int unsigned XLEN = 32,   // is used to quickly switch between 32 and 64 for testing
  // extensions  (see `riscv_isa_pkg` for enumeration definition)
  isa_ext_t    XTEN = RV_M | RV_C | RV_Zicsr,
  // privilige modes
  isa_priv_t   MODES = MODES_M,
  // ISA
  isa_t        ISA = XLEN==32 ? '{spec: '{base: RV_32I , ext: XTEN}, priv: MODES}
                   : XLEN==64 ? '{spec: '{base: RV_64I , ext: XTEN}, priv: MODES}
                              : '{spec: '{base: RV_128I, ext: XTEN}, priv: MODES},
  // instruction bus
  int unsigned IAW = 21,    // instruction address width
  int unsigned IDW = 32,    // instruction data    width
  // data bus
  int unsigned DAW = 17,    // data address width
  int unsigned DDW = XLEN,  // data data    width
  int unsigned DBW = DDW/8  // data byte en width
)(
  // system signals
  input  logic clk,  // clock
  input  logic rst   // reset
);

import riscv_asm_pkg::*;

// clock period counter
int unsigned cnt;
bit timeout = 1'b0;

////////////////////////////////////////////////////////////////////////////////
// DEBUG
////////////////////////////////////////////////////////////////////////////////

initial begin
  $display("==========================================");
  $display("ISA                  : %p", ISA                  );
  $display("ISA.spec             : %b", ISA.spec             );
  $display("ISA.spec.base        : %b", ISA.spec.base        );
  $display("ISA.spec.ext         : %b", ISA.spec.ext         );
  $display("ISA.spec.ext.M       : %b", ISA.spec.ext.M       );
  $display("ISA.spec.ext.A       : %b", ISA.spec.ext.A       );
  $display("ISA.spec.ext.F       : %b", ISA.spec.ext.F       );
  $display("ISA.spec.ext.D       : %b", ISA.spec.ext.D       );
  $display("ISA.spec.ext.Zicsr   : %b", ISA.spec.ext.Zicsr   );
  $display("ISA.spec.ext.Zifencei: %b", ISA.spec.ext.Zifencei);
  $display("ISA.spec.ext.Q       : %b", ISA.spec.ext.Q       );
  $display("ISA.spec.ext.L       : %b", ISA.spec.ext.L       );
  $display("ISA.spec.ext.C       : %b", ISA.spec.ext.C       );
  $display("ISA.spec.ext.B       : %b", ISA.spec.ext.B       );
  $display("ISA.spec.ext.J       : %b", ISA.spec.ext.J       );
  $display("ISA.spec.ext.T       : %b", ISA.spec.ext.T       );
  $display("ISA.spec.ext.P       : %b", ISA.spec.ext.P       );
  $display("ISA.spec.ext.V       : %b", ISA.spec.ext.V       );
  $display("ISA.spec.ext.N       : %b", ISA.spec.ext.N       );
  $display("ISA.spec.ext.H       : %b", ISA.spec.ext.H       );
  $display("ISA.spec.ext.S       : %b", ISA.spec.ext.S       );
  $display("ISA.spec.ext.Zam     : %b", ISA.spec.ext.Zam     );
  $display("ISA.spec.ext.Ztso    : %b", ISA.spec.ext.Ztso    );
  $display("ISA.priv             : %b", ISA.priv             );
  $display("==========================================");
end

////////////////////////////////////////////////////////////////////////////////
// local signals
////////////////////////////////////////////////////////////////////////////////

r5p_bus_if #(.AW (IAW), .DW (IDW)) bus_if (.clk (clk), .rst (rst));
r5p_bus_if #(.AW (DAW), .DW (DDW)) bus_ls (.clk (clk), .rst (rst));

// instruction fetch bus
logic           if_req;
logic [IAW-1:0] if_adr;
logic [IDW-1:0] if_rdt;
logic           if_ack;
// load/store bus, LS memory bus, controller bus
logic           ls_req, ls_mem_req, ls_ctl_req;
logic           ls_wen, ls_mem_wen, ls_ctl_wen;
logic [DAW-1:0] ls_adr, ls_mem_adr, ls_ctl_adr;  // +1 bits for decoder
logic [DBW-1:0] ls_ben, ls_mem_ben, ls_ctl_ben;
logic [DDW-1:0] ls_wdt, ls_mem_wdt, ls_ctl_wdt;
logic [DDW-1:0] ls_rdt, ls_mem_rdt, ls_ctl_rdt;
logic           ls_ack, ls_mem_ack, ls_ctl_ack;

////////////////////////////////////////////////////////////////////////////////
// RTL DUT instance
////////////////////////////////////////////////////////////////////////////////

r5p_core #(
  // RISC-V ISA
  .ISA  (ISA),
  .XLEN (XLEN),
  // instruction bus
  .IDW  (IDW),
  .IAW  (IAW),
  // data bus
  .DAW  (DAW),
  .DDW  (DDW)
) DUT (
  // system signals
  .clk     (clk),
  .rst     (rst),
  // instruction fetch
  .if_req  (bus_if.vld),
  .if_adr  (bus_if.adr),
  .if_rdt  (bus_if.rdt),
  .if_ack  (bus_if.rdy),
  // data load/store
  .ls_req  (bus_ls.vld),
  .ls_wen  (bus_ls.wen),
  .ls_adr  (bus_ls.adr),
  .ls_ben  (bus_ls.ben),
  .ls_wdt  (bus_ls.wdt),
  .ls_rdt  (bus_ls.rdt),
  .ls_ack  (bus_ls.rdy)
);

assign bus_if.wen = 1'b0;
assign bus_if.ben = '1;
assign bus_if.wen = 'x;

////////////////////////////////////////////////////////////////////////////////
// program memory
////////////////////////////////////////////////////////////////////////////////

string if_str;
always if_str = disasm(ISA, if_rdt);

mem #(
  .ISA  (ISA),
  .FN   ("mem_if.bin"),
  .SZ   (2**IAW),
  .DW   (IDW),
  .DBG  ("INS"),
  .OPC  (1'b1)
) mem_if (
  // system signals
  .clk  (clk),
  // instruction fetch
  .req  (bus_if.vld),
  .wen  (bus_if.wen),
  .adr  (bus_if.adr),
  .ben  (bus_if.ben),
  .wdt  (bus_if.wdt),
  .rdt  (bus_if.rdt),
  .ack  (bus_if.rdy)
);

/*
r5p_bus_mon #(
  .DW   (IDW),
  .AW   (IAW),
) bus_mon_if (
  // system signals
  .clk  (clk),
  .rst  (rst),
  // instruction fetch
  .req  (if_req),
  .wen  (1'b0),
  .adr  (if_adr),
  .ben  ('1),
  .wdt  ('x),
  .rdt  (if_rdt),
  .ack  (if_ack)
);
*/

////////////////////////////////////////////////////////////////////////////////
// load/store bus decoder
////////////////////////////////////////////////////////////////////////////////

r5p_bus_dec #(
  .AW  (DAW),
  .DW  (DDW),
  .BN  (2),       // bus number
  .AS  ({ {1'b1, {(DAW-1){1'bx}}} ,   // 0x0_0000 ~ 0x0_ffff - data memory
          {1'b0, {(DAW-1){1'bx}}} })  // 0x1_0000 ~ 0x1_ffff - controller
) ls_dec (
  // system signals
  .clk  (clk),
  .rst  (rst),
  // data load/store
  // slave port and master ports
  .s_req  (bus_ls.vld),  .m_req  ('{ls_ctl_req, ls_mem_req}),
  .s_wen  (bus_ls.wen),  .m_wen  ('{ls_ctl_wen, ls_mem_wen}),
  .s_ben  (bus_ls.ben),  .m_ben  ('{ls_ctl_ben, ls_mem_ben}),
  .s_adr  (bus_ls.adr),  .m_adr  ('{ls_ctl_adr, ls_mem_adr}),
  .s_wdt  (bus_ls.wdt),  .m_wdt  ('{ls_ctl_wdt, ls_mem_wdt}),
  .s_rdt  (bus_ls.rdt),  .m_rdt  ('{ls_ctl_rdt, ls_mem_rdt}),
  .s_ack  (bus_ls.rdy),  .m_ack  ('{ls_ctl_ack, ls_mem_ack})
);

////////////////////////////////////////////////////////////////////////////////
// data memory
////////////////////////////////////////////////////////////////////////////////

mem #(
  .ISA  (ISA),
  .FN   ("mem_ls.bin"),
  .SZ   (2**(DAW-1)),
  .DW   (DDW),
  .DBG  ("DAT"),
  .TXT  (1'b1)
) mem_ls (
  // system signals
  .clk  (clk),
  // data load/store
  .req  (ls_mem_req),
  .wen  (ls_mem_wen),
  .ben  (ls_mem_ben),
  .adr  (ls_mem_adr[DAW-2:0]),
  .wdt  (ls_mem_wdt),
  .rdt  (ls_mem_rdt),
  .ack  (ls_mem_ack)
);

/*
r5p_bus_mon #(
  .DW   (DDW),
  .AW   (DAW),
) bus_mon_ls (
  // system signals
  .clk  (clk),
  .rst  (rst),
  // data load/store
  .req  (ls_req),
  .wen  (ls_wen),
  .adr  (ls_adr),
  .ben  (ls_ben),
  .wdt  (ls_wdt),
  .rdt  (ls_rdt),
  .ack  (ls_ack)
);
*/

////////////////////////////////////////////////////////////////////////////////
// controller
////////////////////////////////////////////////////////////////////////////////

logic [DDW-1:0] rvmodel_data_begin;
logic [DDW-1:0] rvmodel_data_end;
logic           rvmodel_halt = '0;

always_ff @(posedge clk, posedge rst)
if (rst) begin
  rvmodel_data_begin <= 'x;
  rvmodel_data_end   <= 'x;
  rvmodel_halt       <= '0;
end else if (ls_ctl_req & ls_ctl_ack) begin
  if (ls_ctl_wen) begin
    // write access
    case (ls_ctl_adr[5-1:0])
      5'h00:  rvmodel_data_begin <= ls_ctl_wdt;
      5'h08:  rvmodel_data_end   <= ls_ctl_wdt;
      5'h10:  rvmodel_halt       <= ls_ctl_wdt[0];
      default:  ;  // do nothing
    endcase
  end
end

// controller response is immediate
assign ls_ctl_ack = 1'b1;

// finish simulation
always @(posedge clk)
if (rvmodel_halt | timeout) begin
  if (rvmodel_halt)  $display("HALT");
  if (timeout     )  $display("TIMEOUT");
  void'(mem_ls.write_hex("signature_debug.txt", 'h10000200, 'h1000021c));
  void'(mem_ls.write_hex("signature.txt", int'(rvmodel_data_begin), int'(rvmodel_data_end)));
  $finish;
end

// at the end dump the test signature
// TODO: not working in Verilator, at least if the C code ends the simulation.
final begin
  $display("FINAL");
  void'(mem_ls.write_hex("signature.txt", int'(rvmodel_data_begin), int'(rvmodel_data_end)));
  $display("TIME: cnt = %d", cnt);
end

////////////////////////////////////////////////////////////////////////////////
// timeout
////////////////////////////////////////////////////////////////////////////////

// time counter
always_ff @(posedge clk, posedge rst)
if (rst) begin
  cnt <= 0;
end else begin
  cnt <= cnt+1;
end

// timeout
//always @(posedge clk)
//if (cnt > 5000)  timeout <= 1'b1;

////////////////////////////////////////////////////////////////////////////////
// waveforms
////////////////////////////////////////////////////////////////////////////////

//initial begin
//  $dumpfile("rp32_tb.vcd");
//  $dumpvars(0, rp32_tb);
//end

endmodule: r5p_tb