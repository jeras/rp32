package riscv_asm;

typedef struct packed {logic [ 6: 0] func7 ;                                                   logic [ 4: 0] rs2      ; logic [ 4: 0] rs1      ; logic [ 2: 0] func3    ; logic [ 4: 0] rd       ;                       logic [ 6: 0] opcode;} t_format_r ;
typedef struct packed {logic [ 4: 0] rs3   ; logic [ 1: 0] func2    ;                          logic [ 4: 0] rs2      ; logic [ 4: 0] rs1      ; logic [ 2: 0] func3    ; logic [ 4: 0] rd       ;                       logic [ 6: 0] opcode;} t_format_r4;
typedef struct packed {logic [11:11] imm_11; logic [10: 5] imm_10_05; logic [ 4: 1] imm_04_01; logic [ 0: 0] imm_00   ; logic [ 4: 0] rs1      ; logic [ 2: 0] func3    ; logic [ 4: 0] rd       ;                       logic [ 6: 0] opcode;} t_format_i ;
typedef struct packed {logic [11:11] imm_11; logic [10: 5] imm_10_05;                          logic [ 4: 0] rs2      ; logic [ 4: 0] rs1      ; logic [ 2: 0] func3    ; logic [ 4: 1] imm_04_01; logic [ 0: 0] imm_00; logic [ 6: 0] opcode;} t_format_s ;
typedef struct packed {logic [12:12] imm_12; logic [10: 5] imm_10_05;                          logic [ 4: 0] rs2      ; logic [ 4: 0] rs1      ; logic [ 2: 0] func3    ; logic [ 4: 1] imm_04_01; logic [11:11] imm_11; logic [ 6: 0] opcode;} t_format_sb;
typedef struct packed {logic [31:31] imm_31; logic [30:20] imm_30_20; logic [19:15] imm_19_15; logic [14:12] imm_14_12;                                                   logic [ 4: 0] rd       ;                       logic [ 6: 0] opcode;} t_format_u ;
typedef struct packed {logic [20:20] imm_20; logic [10: 5] imm_10_05; logic [ 4: 1] imm_04_01; logic [11:11] imm_11   ; logic [19:15] imm_19_15; logic [14:12] imm_14_12; logic [ 4: 0] rd       ;                       logic [ 6: 0] opcode;} t_format_uj;

typedef union packed {
  t_format_r  r ;
  t_format_r4 r4;
  t_format_i  i ;
  t_format_s  s ;
  t_format_sb sb;
  t_format_u  u ;
  t_format_uj uj;
} t_format;

typedef enum logic [3:0] {TYPE_R, TYPE_R4, TYPE_I, TYPE_L, TYPE_S, TYPE_SB, TYPE_U, TYPE_UJ, TYPE_0, TYPE_X} t_format_sel;

function logic signed [31:0] immediate (t_format i, t_format_sel sel);
  case (sel)
    TYPE_L,
    TYPE_I : immediate = {{21{i.i .imm_11}},                                                              i.i .imm_10_05, i.i .imm_04_01, i.i .imm_00}; // s11
    TYPE_S : immediate = {{21{i.s .imm_11}},                                                              i.s .imm_10_05, i.s .imm_04_01, i.s .imm_00}; // s11
    TYPE_SB: immediate = {{20{i.sb.imm_12}},                                                 i.sb.imm_11, i.sb.imm_10_05, i.sb.imm_04_01, 1'b0       }; // s12
    TYPE_U : immediate = {    i.u .imm_31  , i.u .imm_30_20, i.u .imm_19_15, i.u .imm_14_12, 12'h000                                                 }; // s31
    TYPE_UJ: immediate = {{12{i.uj.imm_20}},                 i.uj.imm_19_15, i.uj.imm_14_12, i.uj.imm_11, i.uj.imm_10_05, i.uj.imm_04_01, 1'b0       }; // s20
    default: immediate = '0; // TODO
  endcase
endfunction: immediate

///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////

typedef struct {
  string               nam;  // name
//  bit [18-1:0] [8-1:0] nam;  // name
  t_format_sel         typ;  // type
//integer              ext;  // extension
} t_asm;

function t_asm decode (t_format opcode);
  casez (opcode)
    //  fedc_ba98_7654_3210_fedc_ba98_7654_3210
    32'b0000_0000_0000_0000_0000_0000_0001_0011: decode = '{"nop               ", TYPE_0 };
    32'b0000_0000_0000_0000_0100_0000_0011_0011: decode = '{"-                 ", TYPE_0 }; // 32'h00004033 - machine generated bubble
    32'b????_????_????_????_?000_????_?110_0011: decode = '{"beq               ", TYPE_SB};
    32'b????_????_????_????_?001_????_?110_0011: decode = '{"bne               ", TYPE_SB};
    32'b????_????_????_????_?100_????_?110_0011: decode = '{"blt               ", TYPE_SB};
    32'b????_????_????_????_?101_????_?110_0011: decode = '{"bge               ", TYPE_SB};
    32'b????_????_????_????_?110_????_?110_0011: decode = '{"bltu              ", TYPE_SB};
    32'b????_????_????_????_?111_????_?110_0011: decode = '{"bgeu              ", TYPE_SB};
    32'b????_????_????_????_?000_????_?110_0111: decode = '{"jalr              ", TYPE_L };
    32'b????_????_????_????_????_????_?110_1111: decode = '{"jal               ", TYPE_UJ};
    32'b????_????_????_????_????_????_?011_0111: decode = '{"lui               ", TYPE_U };
    32'b????_????_????_????_????_????_?001_0111: decode = '{"auipc             ", TYPE_U };
    32'b????_????_????_????_?000_????_?001_0011: decode = '{"addi              ", TYPE_I };
    32'b0000_00??_????_????_?001_????_?001_0011: decode = '{"slli              ", TYPE_R };
    32'b????_????_????_????_?010_????_?001_0011: decode = '{"slti              ", TYPE_I };
    32'b????_????_????_????_?011_????_?001_0011: decode = '{"sltiu             ", TYPE_I };
    32'b????_????_????_????_?100_????_?001_0011: decode = '{"xori              ", TYPE_I };
    32'b0000_00??_????_????_?101_????_?001_0011: decode = '{"srli              ", TYPE_R };
    32'b0100_00??_????_????_?101_????_?001_0011: decode = '{"srai              ", TYPE_R };
    32'b????_????_????_????_?110_????_?001_0011: decode = '{"ori               ", TYPE_I };
    32'b????_????_????_????_?111_????_?001_0011: decode = '{"andi              ", TYPE_I };
    32'b0000_000?_????_????_?000_????_?011_0011: decode = '{"add               ", TYPE_R };
    32'b0100_000?_????_????_?000_????_?011_0011: decode = '{"sub               ", TYPE_R };
    32'b0000_000?_????_????_?001_????_?011_0011: decode = '{"sll               ", TYPE_R };
    32'b0000_000?_????_????_?010_????_?011_0011: decode = '{"slt               ", TYPE_R };
    32'b0000_000?_????_????_?011_????_?011_0011: decode = '{"sltu              ", TYPE_R };
    32'b0000_000?_????_????_?100_????_?011_0011: decode = '{"xor               ", TYPE_R };
    32'b0000_000?_????_????_?101_????_?011_0011: decode = '{"srl               ", TYPE_R };
    32'b0100_000?_????_????_?101_????_?011_0011: decode = '{"sra               ", TYPE_R };
    32'b0000_000?_????_????_?110_????_?011_0011: decode = '{"or                ", TYPE_R };
    32'b0000_000?_????_????_?111_????_?011_0011: decode = '{"and               ", TYPE_R };
    32'b????_????_????_????_?000_????_?001_1011: decode = '{"addiw             ", TYPE_I };
    32'b0000_000?_????_????_?001_????_?001_1011: decode = '{"slliw             ", TYPE_R };
    32'b0000_000?_????_????_?101_????_?001_1011: decode = '{"srliw             ", TYPE_R };
    32'b0100_000?_????_????_?101_????_?001_1011: decode = '{"sraiw             ", TYPE_R };
    32'b0000_000?_????_????_?000_????_?011_1011: decode = '{"addw              ", TYPE_R };
    32'b0100_000?_????_????_?000_????_?011_1011: decode = '{"subw              ", TYPE_R };
    32'b0000_000?_????_????_?001_????_?011_1011: decode = '{"sllw              ", TYPE_R };
    32'b0000_000?_????_????_?101_????_?011_1011: decode = '{"srlw              ", TYPE_R };
    32'b0100_000?_????_????_?101_????_?011_1011: decode = '{"sraw              ", TYPE_R };
    32'b????_????_????_????_?000_????_?000_0011: decode = '{"lb                ", TYPE_L };
    32'b????_????_????_????_?001_????_?000_0011: decode = '{"lh                ", TYPE_L };
    32'b????_????_????_????_?010_????_?000_0011: decode = '{"lw                ", TYPE_L };
    32'b????_????_????_????_?011_????_?000_0011: decode = '{"ld                ", TYPE_L };
    32'b????_????_????_????_?100_????_?000_0011: decode = '{"lbu               ", TYPE_L };
    32'b????_????_????_????_?101_????_?000_0011: decode = '{"lhu               ", TYPE_L };
    32'b????_????_????_????_?110_????_?000_0011: decode = '{"lwu               ", TYPE_L };
    32'b????_????_????_????_?000_????_?010_0011: decode = '{"sb                ", TYPE_S };
    32'b????_????_????_????_?001_????_?010_0011: decode = '{"sh                ", TYPE_S };
    32'b????_????_????_????_?010_????_?010_0011: decode = '{"sw                ", TYPE_S };
    32'b????_????_????_????_?011_????_?010_0011: decode = '{"sd                ", TYPE_S };
    32'b????_????_????_????_?000_????_?000_1111: decode = '{"fence             ", TYPE_0 };
    32'b????_????_????_????_?001_????_?000_1111: decode = '{"fence.i           ", TYPE_0 };
    32'b0000_001?_????_????_?000_????_?011_0011: decode = '{"mul               ", TYPE_R };
    32'b0000_001?_????_????_?001_????_?011_0011: decode = '{"mulh              ", TYPE_R };
    32'b0000_001?_????_????_?010_????_?011_0011: decode = '{"mulhsu            ", TYPE_R };
    32'b0000_001?_????_????_?011_????_?011_0011: decode = '{"mulhu             ", TYPE_R };
    32'b0000_001?_????_????_?100_????_?011_0011: decode = '{"div               ", TYPE_R };
    32'b0000_001?_????_????_?101_????_?011_0011: decode = '{"divu              ", TYPE_R };
    32'b0000_001?_????_????_?110_????_?011_0011: decode = '{"rem               ", TYPE_R };
    32'b0000_001?_????_????_?111_????_?011_0011: decode = '{"remu              ", TYPE_R };
    32'b0000_001?_????_????_?000_????_?011_1011: decode = '{"mulw              ", TYPE_R };
    32'b0000_001?_????_????_?100_????_?011_1011: decode = '{"divw              ", TYPE_R };
    32'b0000_001?_????_????_?101_????_?011_1011: decode = '{"divuw             ", TYPE_R };
    32'b0000_001?_????_????_?110_????_?011_1011: decode = '{"remw              ", TYPE_R };
    32'b0000_001?_????_????_?111_????_?011_1011: decode = '{"remuw             ", TYPE_R };
    32'b0000_0???_????_????_?010_????_?010_1111: decode = '{"amoadd.w          ", TYPE_R };
    32'b0010_0???_????_????_?010_????_?010_1111: decode = '{"amoxor.w          ", TYPE_R };
    32'b0100_0???_????_????_?010_????_?010_1111: decode = '{"amoor.w           ", TYPE_R };
    32'b0110_0???_????_????_?010_????_?010_1111: decode = '{"amoand.w          ", TYPE_R };
    32'b1000_0???_????_????_?010_????_?010_1111: decode = '{"amomin.w          ", TYPE_R };
    32'b1010_0???_????_????_?010_????_?010_1111: decode = '{"amomax.w          ", TYPE_R };
    32'b1100_0???_????_????_?010_????_?010_1111: decode = '{"amominu.w         ", TYPE_R };
    32'b1110_0???_????_????_?010_????_?010_1111: decode = '{"amomaxu.w         ", TYPE_R };
    32'b0000_1???_????_????_?010_????_?010_1111: decode = '{"amoswap.w         ", TYPE_R };
    32'b0001_0??0_0000_????_?010_????_?010_1111: decode = '{"lr.w              ", TYPE_R };
    32'b0001_1???_????_????_?010_????_?010_1111: decode = '{"sc.w              ", TYPE_R };
    32'b0000_0???_????_????_?011_????_?010_1111: decode = '{"amoadd.d          ", TYPE_R };
    32'b0010_0???_????_????_?011_????_?010_1111: decode = '{"amoxor.d          ", TYPE_R };
    32'b0100_0???_????_????_?011_????_?010_1111: decode = '{"amoor.d           ", TYPE_R };
    32'b0110_0???_????_????_?011_????_?010_1111: decode = '{"amoand.d          ", TYPE_R };
    32'b1000_0???_????_????_?011_????_?010_1111: decode = '{"amomin.d          ", TYPE_R };
    32'b1010_0???_????_????_?011_????_?010_1111: decode = '{"amomax.d          ", TYPE_R };
    32'b1100_0???_????_????_?011_????_?010_1111: decode = '{"amominu.d         ", TYPE_R };
    32'b1110_0???_????_????_?011_????_?010_1111: decode = '{"amomaxu.d         ", TYPE_R };
    32'b0000_1???_????_????_?011_????_?010_1111: decode = '{"amoswap.d         ", TYPE_R };
    32'b0001_0??0_0000_????_?011_????_?010_1111: decode = '{"lr.d              ", TYPE_R };
    32'b0001_1???_????_????_?011_????_?010_1111: decode = '{"sc.d              ", TYPE_R };
    32'b0000_0000_0000_0000_0000_0000_0111_0011: decode = '{"scall             ", TYPE_0 };
    32'b0000_0000_0001_0000_0000_0000_0111_0011: decode = '{"sbreak            ", TYPE_0 };
    32'b1000_0000_0000_0000_0000_0000_0111_0011: decode = '{"sret              ", TYPE_0 };
    32'b????_????_????_????_?001_????_?111_0011: decode = '{"csrrw             ", TYPE_I };
    32'b????_????_????_????_?010_????_?111_0011: decode = '{"csrrs             ", TYPE_I };
    32'b????_????_????_????_?011_????_?111_0011: decode = '{"csrrc             ", TYPE_I };
    32'b????_????_????_????_?101_????_?111_0011: decode = '{"csrrwi            ", TYPE_I };
    32'b????_????_????_????_?110_????_?111_0011: decode = '{"csrrsi            ", TYPE_I };
    32'b????_????_????_????_?111_????_?111_0011: decode = '{"csrrci            ", TYPE_I };
    default                                    : decode = '{"csrrci            ", TYPE_X };
  endcase
endfunction: decode

//  '{"fadd_s            ", TYPE_,32'b0000000??????????????????1010011},
//  '{"fsub_s            ", TYPE_,32'b0000100??????????????????1010011},
//  '{"fmul_s            ", TYPE_,32'b0001000??????????????????1010011},
//  '{"fdiv_s            ", TYPE_,32'b0001100??????????????????1010011},
//  '{"fsgnj_s           ", TYPE_,32'b0010000??????????000?????1010011},
//  '{"fsgnjn_s          ", TYPE_,32'b0010000??????????001?????1010011},
//  '{"fsgnjx_s          ", TYPE_,32'b0010000??????????010?????1010011},
//  '{"fmin_s            ", TYPE_,32'b0010100??????????000?????1010011},
//  '{"fmax_s            ", TYPE_,32'b0010100??????????001?????1010011},
//  '{"fsqrt_s           ", TYPE_,32'b010110000000?????????????1010011},
//  '{"fadd_d            ", TYPE_,32'b0000001??????????????????1010011},
//  '{"fsub_d            ", TYPE_,32'b0000101??????????????????1010011},
//  '{"fmul_d            ", TYPE_,32'b0001001??????????????????1010011},
//  '{"fdiv_d            ", TYPE_,32'b0001101??????????????????1010011},
//  '{"fsgnj_d           ", TYPE_,32'b0010001??????????000?????1010011},
//  '{"fsgnjn_d          ", TYPE_,32'b0010001??????????001?????1010011},
//  '{"fsgnjx_d          ", TYPE_,32'b0010001??????????010?????1010011},
//  '{"fmin_d            ", TYPE_,32'b0010101??????????000?????1010011},
//  '{"fmax_d            ", TYPE_,32'b0010101??????????001?????1010011},
//  '{"fcvt_s_d          ", TYPE_,32'b010000000001?????????????1010011},
//  '{"fcvt_d_s          ", TYPE_,32'b010000100000?????????????1010011},
//  '{"fsqrt_d           ", TYPE_,32'b010110100000?????????????1010011},
//  '{"fle_s             ", TYPE_,32'b1010000??????????000?????1010011},
//  '{"flt_s             ", TYPE_,32'b1010000??????????001?????1010011},
//  '{"feq_s             ", TYPE_,32'b1010000??????????010?????1010011},
//  '{"fle_d             ", TYPE_,32'b1010001??????????000?????1010011},
//  '{"flt_d             ", TYPE_,32'b1010001??????????001?????1010011},
//  '{"feq_d             ", TYPE_,32'b1010001??????????010?????1010011},
//  '{"fcvt_w_s          ", TYPE_,32'b110000000000?????????????1010011},
//  '{"fcvt_wu_s         ", TYPE_,32'b110000000001?????????????1010011},
//  '{"fcvt_l_s          ", TYPE_,32'b110000000010?????????????1010011},
//  '{"fcvt_lu_s         ", TYPE_,32'b110000000011?????????????1010011},
//  '{"fmv_x_s           ", TYPE_,32'b111000000000?????000?????1010011},
//  '{"fclass_s          ", TYPE_,32'b111000000000?????001?????1010011},
//  '{"fcvt_w_d          ", TYPE_,32'b110000100000?????????????1010011},
//  '{"fcvt_wu_d         ", TYPE_,32'b110000100001?????????????1010011},
//  '{"fcvt_l_d          ", TYPE_,32'b110000100010?????????????1010011},
//  '{"fcvt_lu_d         ", TYPE_,32'b110000100011?????????????1010011},
//  '{"fmv_x_d           ", TYPE_,32'b111000100000?????000?????1010011},
//  '{"fclass_d          ", TYPE_,32'b111000100000?????001?????1010011},
//  '{"fcvt_s_w          ", TYPE_,32'b110100000000?????????????1010011},
//  '{"fcvt_s_wu         ", TYPE_,32'b110100000001?????????????1010011},
//  '{"fcvt_s_l          ", TYPE_,32'b110100000010?????????????1010011},
//  '{"fcvt_s_lu         ", TYPE_,32'b110100000011?????????????1010011},
//  '{"fmv_s_x           ", TYPE_,32'b111100000000?????000?????1010011},
//  '{"fcvt_d_w          ", TYPE_,32'b110100100000?????????????1010011},
//  '{"fcvt_d_wu         ", TYPE_,32'b110100100001?????????????1010011},
//  '{"fcvt_d_l          ", TYPE_,32'b110100100010?????????????1010011},
//  '{"fcvt_d_lu         ", TYPE_,32'b110100100011?????????????1010011},
//  '{"fmv_d_x           ", TYPE_,32'b111100100000?????000?????1010011},
//  '{"flw               ", TYPE_,32'b?????????????????010?????0000111},
//  '{"fld               ", TYPE_,32'b?????????????????011?????0000111},
//  '{"fsw               ", TYPE_,32'b?????????????????010?????0100111},
//  '{"fsd               ", TYPE_,32'b?????????????????011?????0100111},
//  '{"fmadd_s           ", TYPE_,32'b?????00??????????????????1000011},
//  '{"fmsub_s           ", TYPE_,32'b?????00??????????????????1000111},
//  '{"fnmsub_s          ", TYPE_,32'b?????00??????????????????1001011},
//  '{"fnmadd_s          ", TYPE_,32'b?????00??????????????????1001111},
//  '{"fmadd_d           ", TYPE_,32'b?????01??????????????????1000011},
//  '{"fmsub_d           ", TYPE_,32'b?????01??????????????????1000111},
//  '{"fnmsub_d          ", TYPE_,32'b?????01??????????????????1001011},
//  '{"fnmadd_d          ", TYPE_,32'b?????01??????????????????1001111},
//  '{"custom0           ", TYPE_,32'b?????????????????000?????0001011},
//  '{"custom0_rs1       ", TYPE_,32'b?????????????????010?????0001011},
//  '{"custom0_rs1_rs2   ", TYPE_,32'b?????????????????011?????0001011},
//  '{"custom0_rd        ", TYPE_,32'b?????????????????100?????0001011},
//  '{"custom0_rd_rs1    ", TYPE_,32'b?????????????????110?????0001011},
//  '{"custom0_rd_rs1_rs2", TYPE_,32'b?????????????????111?????0001011},
//  '{"custom1           ", TYPE_,32'b?????????????????000?????0101011},
//  '{"custom1_rs1       ", TYPE_,32'b?????????????????010?????0101011},
//  '{"custom1_rs1_rs2   ", TYPE_,32'b?????????????????011?????0101011},
//  '{"custom1_rd        ", TYPE_,32'b?????????????????100?????0101011},
//  '{"custom1_rd_rs1    ", TYPE_,32'b?????????????????110?????0101011},
//  '{"custom1_rd_rs1_rs2", TYPE_,32'b?????????????????111?????0101011},
//  '{"custom2           ", TYPE_,32'b?????????????????000?????1011011},
//  '{"custom2_rs1       ", TYPE_,32'b?????????????????010?????1011011},
//  '{"custom2_rs1_rs2   ", TYPE_,32'b?????????????????011?????1011011},
//  '{"custom2_rd        ", TYPE_,32'b?????????????????100?????1011011},
//  '{"custom2_rd_rs1    ", TYPE_,32'b?????????????????110?????1011011},
//  '{"custom2_rd_rs1_rs2", TYPE_,32'b?????????????????111?????1011011},
//  '{"custom3           ", TYPE_,32'b?????????????????000?????1111011},
//  '{"custom3_rs1       ", TYPE_,32'b?????????????????010?????1111011},
//  '{"custom3_rs1_rs2   ", TYPE_,32'b?????????????????011?????1111011},
//  '{"custom3_rd        ", TYPE_,32'b?????????????????100?????1111011},
//  '{"custom3_rd_rs1    ", TYPE_,32'b?????????????????110?????1111011},
//  '{"custom3_rd_rs1_rs2", TYPE_,32'b?????????????????111?????1111011},

///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////

parameter string REG_X [0:31] = '{"x0 ", "ra ", "s0 ", "s1 ", "s2 ", "s3 ", "s4 ", "s5 ", "s6 ", "s7 ", "s8 ", "s9 ", "s10", "s11", "sp ", "tp ",
                                  "v0 ", "v1 ", "a0 ", "a1 ", "a2 ", "a3 ", "a4 ", "a5 ", "a6 ", "a7 ", "a8 ", "a9 ", "a10", "a11", "a12", "a13"};
parameter string REG_F [0:31] = '{" fs0"," fs1"," fs2"," fs3"," fs4"," fs5"," fs6"," fs7"," fs8"," fs9","fs10","fs11","fs12","fs13","fs14","fs15",
                                  " fv0"," fv1"," fa0"," fa1"," fa2"," fa3"," fa4"," fa5"," fa6"," fa7"," fa8"," fa9","fa10","fa11","fa12","fa13"};
parameter string REG_P [0:31] = '{" cr0"," cr1"," cr2"," cr3"," cr4"," cr5"," cr6"," cr7"," cr8"," cr9","cr10","cr11","cr12","cr13","cr14","cr15",
                                  "cr16","cr17","cr18","cr19","cr20","cr21","cr22","cr23","cr24","cr25","cr26","cr27","cr28","cr29","cr30","cr31"};

function string reg_x (
  logic [5-1:0] r,
  bit           abi
);
  reg_x = abi ? REG_X[r] : $sformatf("r%0d", r);
endfunction: reg_x

///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////

function string dis (
  t_format code,
  bit      abi=1  // enable "ABI" style register names
);

  logic [32-1:0] imm;
  t_asm op;

  op  = decode(code);
  imm = immediate(code, op.typ);
  case (op.typ)
    TYPE_R :  dis = $sformatf("%s %s, %s, %s"        , op.nam, reg_x(code.r .rd , abi),      reg_x(code.r .rs1, abi), reg_x(code.r .rs2, abi)     );
    TYPE_0 :  dis = $sformatf("%s"                   , op.nam                                                                                     );
    TYPE_I :  dis = $sformatf("%s %s, %s, 0x%03x"    , op.nam, reg_x(code.i .rd , abi),      reg_x(code.i .rs1, abi),                          imm);
    TYPE_SB:  dis = $sformatf("%s %s, %s, 0x%04x"    , op.nam,                               reg_x(code.sb.rs1, abi), reg_x(code.sb.rs2, abi), imm);
    TYPE_UJ:  dis = $sformatf("%s 0x%06x"            , op.nam,                                                                                 imm);
    TYPE_U :  dis = $sformatf("%s %s, 0x%08x"        , op.nam, reg_x(code.u .rd , abi),                                                        imm);
    TYPE_L :  dis = $sformatf("%s %s, 0x%03x (%s)"   , op.nam, reg_x(code.i .rd , abi), imm, reg_x(code.i .rs1, abi),                             );
    TYPE_S :  dis = $sformatf("%s %s, 0x%03x (%s)"   , op.nam, reg_x(code.s .rs2, abi), imm, reg_x(code.s .rs1, abi),                             );
    default:  dis =           "unknown";
  endcase

endfunction

///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////

//function logic [32-1:0] asm (
//  input byte [128-1:0] str;
//);
//endfunction

endpackage: riscv_asm
