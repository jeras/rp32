endpackage: rp_pkg
