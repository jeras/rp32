///////////////////////////////////////////////////////////////////////////////
// RISC-V ISA package
///////////////////////////////////////////////////////////////////////////////

package riscv_isa_pkg;

///////////////////////////////////////////////////////////////////////////////
// ISA base and extensions
// 2-level type `bit` is used for parameters
///////////////////////////////////////////////////////////////////////////////

struct packed {
  // ISA base
  logic e,  // RV32E  - embedded
  logic w,  // RV32I  - word
  logic d,  // RV64I  - double
  logic q   // RV128I - quad
  // extensions
  logic m,  // integer multiplication and division
  logic a,  // atomic
  logic f,  // single-precision floating-point
  logic d,  // double-precision floating-point
  logic q,  // quad-precision floating-point
  logic l,  // decimal precision floating-point
//logic c,  // compressed
  logic b,  // bit manipulation
  logic j,  // dynamically translated languages
  logic t,  // transactional memory
  logic p,  // packed-SIMD
  logic v,  // vector operations
  logic n   // user-level interrupts
} isa_t;

///////////////////////////////////////////////////////////////////////////////
// I base (32E, 32I, 64I, 128I)
// data types
// 4-level type `logic` is used for signals
///////////////////////////////////////////////////////////////////////////////

// generic size type
enum logic [2-1:0] {
  SZ_B = 3'b000;
  SZ_B = 3'b000;
  SZ_H = 3'b001;
  SZ_W = 3'b010;
  SZ_D = 3'b100;
  SZ_Q = 3'b110;
} sz_t;

// PC multiplexer
enum logic [2-1:0] {
  PC_PC2 = 2'b00;  // next   address 32bit instruction
  PC_PC4 = 2'b01;  // next   address 16bit instruction
  PC_ALU = 2'b10;  // branch address
  PC_EPC = 2'b10;  // EPC value from CSR
} pc_t;

// branch type
enum logic [3-1:0] {
  BR_EQ  = 3'b00_0;  //     equal
  BR_NE  = 3'b00_1;  // not equal
  BR_LTS = 3'b10_0;  // less    then            signed
  BR_GES = 3'b10_1;  // greater then or equal   signed
  BR_LTU = 3'b11_0;  // less    then          unsigned
  BR_GEU = 3'b11_1;  // greater then or equal unsigned
  BR_XXX = 3'bxx_x;  // idle
} br_t;

// ALU argument 1 multiplexer (RS1,...)
enum logic {
  A1_GPR = 1'b0;
  A1_PC  = 1'b1;
} a1_t;

// ALU argument 2 multiplexer (RS2,...)
enum logic {
  A2_GPR = 1'b0;
  A2_IMM = 1'b1;
} a2_t;

// ALU operation
enum logic [4-1:0] {
  // adder based instructions
  AO_ADD,  // addition
  AO_SUB,  // subtraction
  AO_LTS,  // less then   signed (not greater then or equal)
  AO_LTU,  // less then unsigned (not greater then or equal)
  // bitwise logical operations
  AO_AND,  // logic AND
  AO_OR ,  // logic OR
  AO_XOR,  // logic XOR
  // barrel shifter
  AO_SLL,  // shift left logical
  AO_SRL,  // shift right logical
  AO_SRA,  // shift right arithmetic
  // copies
  AO_CP1,  // copy rs1
  AO_CP2,  // copy rs2
  // explicit idle
  AO_XXX,  // do nothing
} alu_t;

// ALU result width
enum logic [2-1:0] {
  AR_S = 2'b00;  // XW
  AR_W = 2'b01;  // word
  AR_D = 2'b10;  // double
  AR_Q = 2'b11;  // quad
} ar_t;

// TODO: check AXI4 encoding for transfer size

// store type
enum logic [3-1:0] {
  ST_B = SZ_B;
  ST_H = SZ_H;
  ST_W = SZ_W;
  ST_D = SZ_D;
  ST_Q = SZ_Q;
} st_t;

// load type
enum logic [4-1:0] {
  LD_B  = {1'b0, SZ_B};  LD_BU = {1'b1, SZ_B};
  LD_H  = {1'b0, SZ_H};  LD_HU = {1'b1, SZ_H};
  LD_W  = {1'b0, SZ_W};  LD_WU = {1'b1, SZ_W};
  LD_D  = {1'b0, SZ_D};  LD_DU = {1'b1, SZ_D};
  LD_Q  = {1'b0, SZ_Q};  LD_QU = {1'b1, SZ_Q};
} ld_t;

// write back multiplexer
enum logic [3-1:0] {
  WB_ALU = 2'b00;
  WB_MEM = 2'b01;
  WB_PC4 = 2'b10;
  WB_CSR = 2'b11;
} wb_t;

// control structure
typedef struct packed {
  pc_t   pc,   // PC multiplexer
  br_t   br,   // branch type
  a1_t   a1,   // ALU RS1 multiplexer
  a2_t   a2,  // ALU RS1 multiplexer
  frm32_t   imm,  // immediate select
  alu_t  alu,  // ALU operation
  sz_t   sza,  // ALU operation size
  st_t   st,   // store type
  logic  ste,  // store enable
  ld_t   ld,   // load type
  logic  lde,  // load enable
  wb_t   wb,   // write back multiplexer
  logic  wbe,  // write back enable
  logic  csr,  // CSR operation
  logic  ill   // illegal
} ctli_t;

///////////////////////////////////////////////////////////////////////////////
// M extension
///////////////////////////////////////////////////////////////////////////////

// M operation
enum logic [2-1:0] {
  MOP_MUL = 2'b00;  // multiplication lower  half result
  MOP_MUH = 2'b01;  // multiplication higher half result
  MOP_DIV = 2'b10;  // division
  MOP_REM = 2'b11;  // reminder
} mop_t;

// control structure
typedef struct packed {
  mop_t op,  // operation
  logic s1,  // sign operand 1
  logic s2,  // sign operand 2
  logic xw,  // XWIDTH (0 - full width, 1 - M64 additional opcodes)
  logic en   // enable
} ctlm_t;


// RV.A32
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                 pc,     rs1,     rs2,   imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b0001_0??0_0000_????_?010_????_?010_1111}: dec32 = '{"lr.w              ", TYPE_32_R};
{16'b????_????????????, 32'b0001_1???_????_????_?010_????_?010_1111}: dec32 = '{"sc.w              ", TYPE_32_R};
{16'b????_????????????, 32'b0000_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoadd.w          ", TYPE_32_R};
{16'b????_????????????, 32'b0010_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoxor.w          ", TYPE_32_R};
{16'b????_????????????, 32'b0100_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoor.w           ", TYPE_32_R};
{16'b????_????????????, 32'b0110_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoand.w          ", TYPE_32_R};
{16'b????_????????????, 32'b1000_0???_????_????_?010_????_?010_1111}: dec32 = '{"amomin.w          ", TYPE_32_R};
{16'b????_????????????, 32'b1010_0???_????_????_?010_????_?010_1111}: dec32 = '{"amomax.w          ", TYPE_32_R};
{16'b????_????????????, 32'b1100_0???_????_????_?010_????_?010_1111}: dec32 = '{"amominu.w         ", TYPE_32_R};
{16'b????_????????????, 32'b1110_0???_????_????_?010_????_?010_1111}: dec32 = '{"amomaxu.w         ", TYPE_32_R};
{16'b????_????????????, 32'b0000_1???_????_????_?010_????_?010_1111}: dec32 = '{"amoswap.w         ", TYPE_32_R};

// RV.A64
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                 pc,     rs1,     rs2,   imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b0001_0??0_0000_????_?011_????_?010_1111}: dec32 = '{"lr.d              ", TYPE_32_R};
{16'b????_????????????, 32'b0001_1???_????_????_?011_????_?010_1111}: dec32 = '{"sc.d              ", TYPE_32_R};
{16'b????_????????????, 32'b0000_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoadd.d          ", TYPE_32_R};
{16'b????_????????????, 32'b0010_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoxor.d          ", TYPE_32_R};
{16'b????_????????????, 32'b0100_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoor.d           ", TYPE_32_R};
{16'b????_????????????, 32'b0110_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoand.d          ", TYPE_32_R};
{16'b????_????????????, 32'b1000_0???_????_????_?011_????_?010_1111}: dec32 = '{"amomin.d          ", TYPE_32_R};
{16'b????_????????????, 32'b1010_0???_????_????_?011_????_?010_1111}: dec32 = '{"amomax.d          ", TYPE_32_R};
{16'b????_????????????, 32'b1100_0???_????_????_?011_????_?010_1111}: dec32 = '{"amominu.d         ", TYPE_32_R};
{16'b????_????????????, 32'b1110_0???_????_????_?011_????_?010_1111}: dec32 = '{"amomaxu.d         ", TYPE_32_R};
{16'b????_????????????, 32'b0000_1???_????_????_?011_????_?010_1111}: dec32 = '{"amoswap.d         ", TYPE_32_R};

///////////////////////////////////////////////////////////////////////////////
// full control structure
///////////////////////////////////////////////////////////////////////////////

// control structure
typedef struct packed {
  ctli_t  i,  // integer
  ctlm_t  m,  // integer multiplication and division
  ctla_t  a,  // atomic
  ctlf_t  f,  // single-precision floating-point
  ctld_t  d,  // double-precision floating-point
  ctlq_t  q,  // quad-precision floating-point
  ctll_t  l,  // decimal precision floating-point
  ctlb_t  b,  // bit manipulation
  ctlj_t  j,  // dynamically translated languages
  ctlt_t  t,  // transactional memory
  ctlp_t  p,  // packed-SIMD
  ctlv_t  v,  // vector operations
  ctln_t  n   // user-level interrupts
} ctl_t;

///////////////////////////////////////////////////////////////////////////////
// instruction size
///////////////////////////////////////////////////////////////////////////////

function int unsigned opsiz (logic [16-1:0] op);
       if (op =?= 16'bx111_xxxx_x111_111)  opsiz = 192;
  else if (op =?= 16'bxxxx_xxxx_x1111111)  opsiz = 80 + 16 * op[14:12];
  else if (op =?= 16'bxxxx_xxxx_x0111111)  opsiz = 64;
  else if (op =?= 16'bxxxx_xxxx_xx011111)  opsiz = 48;
  else if (op !?= 16'bxxxx_xxxx_xxx111xx
       &&  op =?= 16'bxxxx_xxxx_xxxxxx11)  opsiz = 32;
  else                                     opsiz = 16;
endfunction: opsiz

///////////////////////////////////////////////////////////////////////////////
// 32 bit instruction format
///////////////////////////////////////////////////////////////////////////////

typedef struct packed {logic [4:0] rs3; logic [1:0] func2;          logic [4:0] rs2; logic [4:0] rs1; logic [2:0] func3; logic [4:0] rd     ;                       logic [6:0] opcode;} frm_r4;
typedef struct packed {                 logic [6:0] func7;          logic [4:0] rs2; logic [4:0] rs1; logic [2:0] func3; logic [4:0] rd     ;                       logic [6:0] opcode;} frm_r;
typedef struct packed {logic [11:00] imm_11_0;                                       logic [4:0] rs1; logic [2:0] func3; logic [4:0] rd     ;                       logic [6:0] opcode;} frm_i;
typedef struct packed {logic [11:05] imm_11_5;                      logic [4:0] rs2; logic [4:0] rs1; logic [2:0] func3; logic [4:0] imm_4_0;                       logic [6:0] opcode;} frm_s;
typedef struct packed {logic [12:12] imm_12; logic [10:5] imm_10_5; logic [4:0] rs2; logic [4:0] rs1; logic [2:0] func3; logic [4:1] imm_4_1; logic [11:11] imm_11; logic [6:0] opcode;} frm_b;
typedef struct packed {logic [31:12] imm_31_12;                                                                          logic [4:0] rd     ;                       logic [6:0] opcode;} frm_u;
typedef struct packed {logic [20:20] imm_20; logic [10:1] imm_10_1; logic [11:11] imm_11; logic [19:12] imm_19_12;       logic [4:0] rd     ;                       logic [6:0] opcode;} frm_j;

typedef union packed {
  frm_r4 r4;
  frm_r r;
  frm_i i;
  frm_s s;
  frm_b b;
  frm_u u;
  frm_j j;
} frm32_t;

typedef enum logic [3:0] {
  T32_R4,
  T32_R,
  T32_I,
  T32_S,
  T32_B,
  T32_U,
  T32_J
} frm_sel_t;

function logic signed [32-1:0] imm32 (t_format_32 i, t_format_sel sel);
  case (sel)
    T32_R4,
    T32_R: imm32 = 'x;
    T32_I: imm32 = {{20{i[31]}},        i[30:25], i[24:21], i[20]}; // s11
    T32_S: imm32 = {{20{i[31]}},        i[30:25], i[11:08], i[07]}; // s11
    T32_B: imm32 = {{19{i[31]}}, i[07], i[30:25], i[11:08], 1'b0 }; // s12
    T32_U: imm32 = {    i[31:12], 12'h000}; // s31
    T32_J: imm32 = {{12{i[31]}}, i[19:12], i[20], i[30:25], i[24:21], 1'b0}; // s20
    default:   imm32 = 'x;
  endcase
endfunction: imm32

function ctli_t dec32 (isa_t isa, frm32_t op);
// default values
//              pc,    rs1,    rs2,  imm,     alu,   ar,    br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
dec32.i = '{PC_PC4, A1_RS1, A2_RS2,   'x,      'x,   'x,    'x,   'x, '0,    'x, '0,     'x, '0,    'x, '0};
//         {op, s1, s2, xw, en}
dec32.m = '{'x, 'x, 'x, 'x, '0};

casez ({isa, ext, op})
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                   pc,    rs1,    rs2,  imm,     alu,   ar,    br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b0000_0000_0000_0000_0000_0000_0001_0011}: dec32.i = '{PC_PC4,     'x,     'x,   'x,      'x,   'x,    'x,   'x, '0,    'x, '0,     'x, '0,    'x, '0}; // 32'000000013 - nop
{16'b????_????????????, 32'b0000_0000_0000_0000_0100_0000_0011_0011}: dec32.i = '{PC_PC4,     'x,     'x,   'x,      'x,   'x,    'x,   'x, '0,    'x, '0,     'x, '0,    'x, '0}; // 32'h00004033 - machine gen. bubble

// RV.I32
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                   pc,    rs1,    rs2,  imm,     alu,   ar,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b????_????_????_????_????_????_?011_0111}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_U, AO_CPB,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // lui
{16'b????_????????????, 32'b????_????_????_????_????_????_?001_0111}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_U, AO_ADD, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // auipc
{16'b????_????????????, 32'b????_????_????_????_????_????_?110_1111}: dec32.i = '{PC_ALU, A1_PC , A2_IMM, IMM_J, AO_ADD, AR_X,     'x,   'x, '0,    'x, '0, WB_PC4, '1, CSR_N, '0};  // jal
{16'b????_????????????, 32'b????_????_????_????_?000_????_?110_0111}: dec32.i = '{PC_ALU, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0,    'x, '0, WB_PC4, '1, CSR_N, '0};  // jalr
{16'b????_????????????, 32'b????_????_????_????_?000_????_?110_0011}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_B, AO_ADD, AR_X, BR_EQ ,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // beq
{16'b????_????????????, 32'b????_????_????_????_?001_????_?110_0011}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_B, AO_ADD, AR_X, BR_NE ,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // bne
{16'b????_????????????, 32'b????_????_????_????_?100_????_?110_0011}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_B, AO_ADD, AR_X, BR_LT ,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // blt
{16'b????_????????????, 32'b????_????_????_????_?101_????_?110_0011}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_B, AO_ADD, AR_X, BR_GE ,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // bge
{16'b????_????????????, 32'b????_????_????_????_?110_????_?110_0011}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_B, AO_ADD, AR_X, BR_LTU,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // bltu
{16'b????_????????????, 32'b????_????_????_????_?111_????_?110_0011}: dec32.i = '{PC_PC4, A1_PC , A2_IMM, IMM_B, AO_ADD, AR_X, BR_GEU,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // bgeu
{16'b????_????????????, 32'b????_????_????_????_?000_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_B , '1, WB_MEM, '1, CSR_N, '0};  // lb
{16'b????_????????????, 32'b????_????_????_????_?001_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_H , '1, WB_MEM, '1, CSR_N, '0};  // lh
{16'b????_????????????, 32'b????_????_????_????_?010_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_W , '1, WB_MEM, '1, CSR_N, '0};  // lw
{16'b????_????????????, 32'b????_????_????_????_?100_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_BU, '1, WB_MEM, '1, CSR_N, '0};  // lbu
{16'b????_????????????, 32'b????_????_????_????_?101_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_HU, '1, WB_MEM, '1, CSR_N, '0};  // lhu
{16'b????_????????????, 32'b????_????_????_????_?000_????_?010_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_S, AO_ADD, AR_X,     'x, ST_B, '1,    'x, '0,     'x, '0, CSR_N, '0};  // sb
{16'b????_????????????, 32'b????_????_????_????_?001_????_?010_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_S, AO_ADD, AR_X,     'x, ST_H, '1,    'x, '0,     'x, '0, CSR_N, '0};  // sh
{16'b????_????????????, 32'b????_????_????_????_?010_????_?010_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_S, AO_ADD, AR_X,     'x, ST_W, '1,    'x, '0,     'x, '0, CSR_N, '0};  // sw
{16'b????_????????????, 32'b????_????_????_????_?000_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // addi
{16'b????_????????????, 32'b????_????_????_????_?010_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_LTS,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // slti
{16'b????_????????????, 32'b????_????_????_????_?011_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_LTU,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sltiu
{16'b????_????????????, 32'b????_????_????_????_?100_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_XOR,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // xori
{16'b????_????????????, 32'b????_????_????_????_?110_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_OR ,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // ori
{16'b????_????????????, 32'b????_????_????_????_?111_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_AND,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // andi
{16'b????_????????????, 32'b0000_000?_????_????_?001_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SLL, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, |imm[6:$clog2(xw)]};  // slli
{16'b????_????????????, 32'b0000_000?_????_????_?101_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SRL, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, |imm[6:$clog2(xw)]};  // srli
{16'b????_????????????, 32'b0100_000?_????_????_?101_????_?001_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SRA, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, |imm[6:$clog2(xw)]};  // srai
{16'b????_????????????, 32'b0000_000?_????_????_?000_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_ADD, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // add
{16'b????_????????????, 32'b0100_000?_????_????_?000_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SUB, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sub
{16'b????_????????????, 32'b0000_000?_????_????_?010_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_LTS,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // slt
{16'b????_????????????, 32'b0000_000?_????_????_?011_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_LTU,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sltu
{16'b????_????????????, 32'b0000_000?_????_????_?100_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_XOR,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // xor
{16'b????_????????????, 32'b0000_000?_????_????_?001_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SLL, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sll
{16'b????_????????????, 32'b0000_000?_????_????_?101_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SRL, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // srl
{16'b????_????????????, 32'b0100_000?_????_????_?101_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SRA, AR_X,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sra
{16'b????_????????????, 32'b0000_000?_????_????_?110_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_OR ,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // or
{16'b????_????????????, 32'b0000_000?_????_????_?111_????_?011_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_AND,   'x,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // and
{16'b????_????????????, 32'b????_????_????_????_?000_????_?000_1111}: dec32.i = '{PC_PC4,     'x,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // fence
{16'b????_????????????, 32'b????_????_????_????_?001_????_?000_1111}: dec32.i = '{PC_PC4,     'x,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // fence.i
{16'b????_????????????, 32'b????_????_????_????_?001_????_?111_0011}: dec32.i = '{PC_PC4, A1_RS1,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0, WB_CSR, '1, CSR_W, '0};  // csrrw
{16'b????_????????????, 32'b????_????_????_????_?010_????_?111_0011}: dec32.i = '{PC_PC4, A1_RS1,     'x,    'x, AO_CP1,   'x,     'x,   'x, '0,    'x, '0, WB_CSR, '1, CSR_S, '0};  // csrrs
{16'b????_????????????, 32'b????_????_????_????_?011_????_?111_0011}: dec32.i = '{PC_PC4, A1_RS1,     'x,    'x, AO_CP1,   'x,     'x,   'x, '0,    'x, '0, WB_CSR, '1, CSR_C, '0};  // csrrc
{16'b????_????????????, 32'b????_????_????_????_?101_????_?111_0011}: dec32.i = '{PC_PC4,     'x,     'x, IMM_Z,     'x,   'x,     'x,   'x, '0,    'x, '0, WB_CSR, '1, CSR_W, '0};  // csrrwi
{16'b????_????????????, 32'b????_????_????_????_?110_????_?111_0011}: dec32.i = '{PC_PC4,     'x,     'x, IMM_Z,     'x,   'x,     'x,   'x, '0,    'x, '0, WB_CSR, '1, CSR_S, '0};  // csrrsi
{16'b????_????????????, 32'b????_????_????_????_?111_????_?111_0011}: dec32.i = '{PC_PC4,     'x,     'x, IMM_Z,     'x,   'x,     'x,   'x, '0,    'x, '0, WB_CSR, '1, CSR_C, '0};  // csrrci
{16'b????_????????????, 32'b0000_0000_0000_0000_0000_0000_0111_0011}: dec32.i = '{PC_PC4,     'x,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0,     'x, '0, CSR_P, '0};  // ecall
{16'b????_????????????, 32'b0000_0000_0001_0000_0000_0000_0111_0011}: dec32.i = '{PC_PC4,     'x,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0,     'x, '0, CSR_P, '0};  // ebreak
{16'b????_????????????, 32'b0001_0000_0000_0000_0000_0000_0111_0011}: dec32.i = '{PC_EPC,     'x,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0,     'x, '0, CSR_P, '0};  // eret
{16'b????_????????????, 32'b0001_0000_0010_0000_0000_0000_0111_0011}: dec32.i = '{PC_PC4,     'x,     'x,    'x,     'x,   'x,     'x,   'x, '0,    'x, '0,     'x, '0, CSR_N, '0};  // wfi

// RV.I64
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                   pc,    rs1,    rs2,   imm,    alu,   ar,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b00??_????????????, 32'b????_????_????_????_?011_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_D , '1, WB_MEM, '1, CSR_N, '0};  // ld
{16'b00??_????????????, 32'b????_????_????_????_?110_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_WU, '1, WB_MEM, '1, CSR_N, '0};  // lwu
{16'b00??_????????????, 32'b????_????_????_????_?011_????_?010_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_S, AO_ADD, AR_X,     'x, ST_D, '1,    'x, '0,     'x, '0, CSR_N, '0};  // sd
{16'b00??_????????????, 32'b????_????_????_????_?000_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // addiw
{16'b00??_????????????, 32'b0000_000?_????_????_?001_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SLL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, |imm[6:$clog2(xw)]};  // slliw
{16'b00??_????????????, 32'b0000_000?_????_????_?101_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SRL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, |imm[6:$clog2(xw)]};  // srliw
{16'b00??_????????????, 32'b0100_000?_????_????_?101_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SRA, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, |imm[6:$clog2(xw)]};  // sraiw
{16'b00??_????????????, 32'b0000_000?_????_????_?000_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_ADD, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // addw
{16'b00??_????????????, 32'b0100_000?_????_????_?000_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SUB, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // subw
{16'b00??_????????????, 32'b0000_000?_????_????_?001_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SLL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sllw
{16'b00??_????????????, 32'b0000_000?_????_????_?101_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SRL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // srlw
{16'b00??_????????????, 32'b0100_000?_????_????_?101_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SRA, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sraw

// RV.I128
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                   pc,    rs1,    rs2,   imm,    alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b0??1_????????????, 32'b????_????_????_????_?011_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_D , '1, WB_MEM, '1, CSR_N, '0};  // lq
{16'b0??1_????????????, 32'b????_????_????_????_?110_????_?000_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_X,     'x,   'x, '0, LD_WU, '1, WB_MEM, '1, CSR_N, '0};  // ldu
{16'b0??1_????????????, 32'b????_????_????_????_?011_????_?010_0011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_S, AO_ADD, AR_X,     'x, ST_D, '1,    'x, '0,     'x, '0, CSR_N, '0};  // sq
{16'b0??1_????????????, 32'b????_????_????_????_?000_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_ADD, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // addiw
{16'b0??1_????????????, 32'b0000_000?_????_????_?001_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SLL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '???};  // slliw
{16'b0??1_????????????, 32'b0000_000?_????_????_?101_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SRL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '???};  // srliw
{16'b0??1_????????????, 32'b0100_000?_????_????_?101_????_?001_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_IMM, IMM_I, AO_SRA, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '???};  // sraiw
{16'b0??1_????????????, 32'b0000_000?_????_????_?000_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_ADD, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // addw
{16'b0??1_????????????, 32'b0100_000?_????_????_?000_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SUB, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // subw
{16'b0??1_????????????, 32'b0000_000?_????_????_?001_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SLL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sllw
{16'b0??1_????????????, 32'b0000_000?_????_????_?101_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SRL, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // srlw
{16'b0??1_????????????, 32'b0100_000?_????_????_?101_????_?011_1011}: dec32.i = '{PC_PC4, A1_RS1, A2_RS2,    'x, AO_SRA, AR_W,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // sraw

// RV.M32
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210              {     op, s1, s2, xw, en}
{16'b????_1???????????, 32'b0000_001?_????_????_?000_????_?011_0011}: dec32.m = '{MOP_MUL, '1, '1, '0, '1};  // mul
{16'b????_1???????????, 32'b0000_001?_????_????_?001_????_?011_0011}: dec32.m = '{MOP_MUH, '1, '1, '0, '1};  // mulh
{16'b????_1???????????, 32'b0000_001?_????_????_?010_????_?011_0011}: dec32.m = '{MOP_MUH, '1, '0, '0, '1};  // mulhsu
{16'b????_1???????????, 32'b0000_001?_????_????_?011_????_?011_0011}: dec32.m = '{MOP_MUH, '0, '0, '0, '1};  // mulhu
{16'b????_1???????????, 32'b0000_001?_????_????_?100_????_?011_0011}: dec32.m = '{MOP_DIV, '1, '1, '0, '1};  // div
{16'b????_1???????????, 32'b0000_001?_????_????_?101_????_?011_0011}: dec32.m = '{MOP_DIV, '1, '0, '0, '1};  // divu
{16'b????_1???????????, 32'b0000_001?_????_????_?110_????_?011_0011}: dec32.m = '{MOP_REM, '1, '1, '0, '1};  // rem
{16'b????_1???????????, 32'b0000_001?_????_????_?111_????_?011_0011}: dec32.m = '{MOP_REM, '1, '0, '0, '1};  // remu

// RV.M64
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210              {     op, s1, s2, xw, en}
{16'b00??_1???????????, 32'b0000_001?_????_????_?000_????_?011_1011}: dec32.m = '{MOP_MUL, '1, '1, '1, '1};  // mulw
{16'b00??_1???????????, 32'b0000_001?_????_????_?100_????_?011_1011}: dec32.m = '{MOP_DIV, '1, '1, '1, '1};  // divw
{16'b00??_1???????????, 32'b0000_001?_????_????_?101_????_?011_1011}: dec32.m = '{MOP_DIV, '1, '0, '1, '1};  // divuw
{16'b00??_1???????????, 32'b0000_001?_????_????_?110_????_?011_1011}: dec32.m = '{MOP_REM, '1, '1, '1, '1};  // remw
{16'b00??_1???????????, 32'b0000_001?_????_????_?111_????_?011_1011}: dec32.m = '{MOP_REM, '1, '0, '1, '1};  // remuw

// RV.A32
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                 pc,     rs1,     rs2,   imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b0001_0??0_0000_????_?010_????_?010_1111}: dec32 = '{"lr.w              ", TYPE_32_R};
{16'b????_????????????, 32'b0001_1???_????_????_?010_????_?010_1111}: dec32 = '{"sc.w              ", TYPE_32_R};
{16'b????_????????????, 32'b0000_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoadd.w          ", TYPE_32_R};
{16'b????_????????????, 32'b0010_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoxor.w          ", TYPE_32_R};
{16'b????_????????????, 32'b0100_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoor.w           ", TYPE_32_R};
{16'b????_????????????, 32'b0110_0???_????_????_?010_????_?010_1111}: dec32 = '{"amoand.w          ", TYPE_32_R};
{16'b????_????????????, 32'b1000_0???_????_????_?010_????_?010_1111}: dec32 = '{"amomin.w          ", TYPE_32_R};
{16'b????_????????????, 32'b1010_0???_????_????_?010_????_?010_1111}: dec32 = '{"amomax.w          ", TYPE_32_R};
{16'b????_????????????, 32'b1100_0???_????_????_?010_????_?010_1111}: dec32 = '{"amominu.w         ", TYPE_32_R};
{16'b????_????????????, 32'b1110_0???_????_????_?010_????_?010_1111}: dec32 = '{"amomaxu.w         ", TYPE_32_R};
{16'b????_????????????, 32'b0000_1???_????_????_?010_????_?010_1111}: dec32 = '{"amoswap.w         ", TYPE_32_R};

// RV.A64
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                 pc,     rs1,     rs2,   imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b0001_0??0_0000_????_?011_????_?010_1111}: dec32 = '{"lr.d              ", TYPE_32_R};
{16'b????_????????????, 32'b0001_1???_????_????_?011_????_?010_1111}: dec32 = '{"sc.d              ", TYPE_32_R};
{16'b????_????????????, 32'b0000_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoadd.d          ", TYPE_32_R};
{16'b????_????????????, 32'b0010_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoxor.d          ", TYPE_32_R};
{16'b????_????????????, 32'b0100_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoor.d           ", TYPE_32_R};
{16'b????_????????????, 32'b0110_0???_????_????_?011_????_?010_1111}: dec32 = '{"amoand.d          ", TYPE_32_R};
{16'b????_????????????, 32'b1000_0???_????_????_?011_????_?010_1111}: dec32 = '{"amomin.d          ", TYPE_32_R};
{16'b????_????????????, 32'b1010_0???_????_????_?011_????_?010_1111}: dec32 = '{"amomax.d          ", TYPE_32_R};
{16'b????_????????????, 32'b1100_0???_????_????_?011_????_?010_1111}: dec32 = '{"amominu.d         ", TYPE_32_R};
{16'b????_????????????, 32'b1110_0???_????_????_?011_????_?010_1111}: dec32 = '{"amomaxu.d         ", TYPE_32_R};
{16'b????_????????????, 32'b0000_1???_????_????_?011_????_?010_1111}: dec32 = '{"amoswap.d         ", TYPE_32_R};

// RV.F32
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                 pc,     rs1,     rs2,   imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
{16'b????_????????????, 32'b????_????_????_????_?010_????_?000_0111}: dec32 = '{"flw               ", TYPE_32_I};
{16'b????_????????????, 32'b????_????_????_????_?010_????_?010_0111}: dec32 = '{"fsw               ", TYPE_32_S};
{16'b????_????????????, 32'b????_?00?_????_????_????_????_?100_0011}: dec32 = '{"fmadd.s           ", TYPE_32_R4};
{16'b????_????????????, 32'b????_?00?_????_????_????_????_?100_0111}: dec32 = '{"fmsub.s           ", TYPE_32_R4};
{16'b????_????????????, 32'b????_?00?_????_????_????_????_?100_1011}: dec32 = '{"fnmsub.s          ", TYPE_32_R4};
{16'b????_????????????, 32'b????_?00?_????_????_????_????_?100_1111}: dec32 = '{"fnmadd.s          ", TYPE_32_R4};
{16'b????_????????????, 32'b0000_000?_????_????_????_????_?101_0011}: dec32 = '{"fadd.s            ", TYPE_32_R};
{16'b????_????????????, 32'b0000_100?_????_????_????_????_?101_0011}: dec32 = '{"fsub.s            ", TYPE_32_R};
{16'b????_????????????, 32'b0001_000?_????_????_????_????_?101_0011}: dec32 = '{"fmul.s            ", TYPE_32_R};
{16'b????_????????????, 32'b0001_100?_????_????_????_????_?101_0011}: dec32 = '{"fdiv.s            ", TYPE_32_R};
{16'b????_????????????, 32'b0101_1000_0000_????_????_????_?101_0011}: dec32 = '{"fsqrt.s           ", TYPE_32_R};
{16'b????_????????????, 32'b0010_000?_????_????_?000_????_?101_0011}: dec32 = '{"fsgnj.s           ", TYPE_32_R};
{16'b????_????????????, 32'b0010_000?_????_????_?001_????_?101_0011}: dec32 = '{"fsgnjn.s          ", TYPE_32_R};
{16'b????_????????????, 32'b0010_000?_????_????_?010_????_?101_0011}: dec32 = '{"fsgnjx.s          ", TYPE_32_R};
{16'b????_????????????, 32'b0010_100?_????_????_?000_????_?101_0011}: dec32 = '{"fmin.s            ", TYPE_32_R};
{16'b????_????????????, 32'b0010_100?_????_????_?001_????_?101_0011}: dec32 = '{"fmax.s            ", TYPE_32_R};
{16'b????_????????????, 32'b1100_0000_0000_????_????_????_?101_0011}: dec32 = '{"fcvt.w.s          ", TYPE_32_R};
{16'b????_????????????, 32'b1100_0000_0001_????_????_????_?101_0011}: dec32 = '{"fcvt.wu.s         ", TYPE_32_R};
{16'b????_????????????, 32'b1110_0000_0000_????_????_????_?101_0011}: dec32 = '{"fmv.x.w           ", TYPE_32_R};

{16'b????_????????????, 32'b0001_0??0_0000_????_?011_????_?010_1111}: dec32 = '{"lr.d              ", TYPE_32_R};

// RV.F64
//   ewdq mafdqlbjtpvn      fedc_ba98_7654_3210_fedc_ba98_7654_3210                 pc,     rs1,     rs2,   imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill


// 32'b1000_0000_0000_0000_0000_0000_0111_0011: dec32 = '{"sret              ", TYPE_32_0};
default                                                               dec32 = '{PC_PC4,     'x,     'x,   'x,      'x,   'x,    'x,   'x, '0,    'x, '0,     'x, '0,    'x, '0}; // 32'000000013 - nop
endcase
endfunction: dec32

///////////////////////////////////////////////////////////////////////////////
// 16 bit instruction format
///////////////////////////////////////////////////////////////////////////////

typedef struct packed {logic [ 3: 0] funct4;                          logic [ 4: 0] rd_rs1;                          logic [ 4: 0] rs2 ; logic [1:0] opcode;} frm_cr;
typedef struct packed {logic [ 2: 0] funct3; logic [12:12] imm_12_12; logic [ 4: 0] rd_rs1; logic [ 6: 2] imm_06_02;                     logic [1:0] opcode;} frm_ci;
typedef struct packed {logic [ 2: 0] funct3; logic [12: 7] imm_12_07; logic [ 4: 0] rd_rs1;                          logic [ 4: 0] rs2 ; logic [1:0] opcode;} frm_css;
typedef struct packed {logic [ 2: 0] funct3; logic [12: 5] imm_12_05;                                                logic [ 2: 0] rd_ ; logic [1:0] opcode;} frm_ciw;
typedef struct packed {logic [ 2: 0] funct3; logic [12:10] imm_12_10; logic [ 2: 0] rs1_  ; logic [ 6: 5] imm_06_05; logic [ 2: 0] rd_ ; logic [1:0] opcode;} frm_cl;
typedef struct packed {logic [ 2: 0] funct3; logic [12:10] imm_12_10; logic [ 2: 0] rs1_  ; logic [ 6: 5] imm_06_05; logic [ 2: 0] rs2_; logic [1:0] opcode;} frm_cs;
typedef struct packed {logic [ 2: 0] funct3; logic [12:10] off_12_10; logic [ 2: 0] rs1_  ; logic [ 6: 2] off_06_02;                     logic [1:0] opcode;} frm_cb;
typedef struct packed {logic [ 2: 0] funct3; logic [12: 2] target;                                                                       logic [1:0] opcode;} frm_cj;

typedef union packed {
  frm_cr  cr;
  frm_ci  ci;
  frm_css css;
  frm_ciw ciw;
  frm_cl  cl;
  frm_cs  cs;
  frm_cb  cb;
  frm_cj  cj;
} t_format_16;

typedef enum logic [3:0] {
  T16_CR,
  T16_CI,
  T16_CSS,
  T16_CIW,
  T16_CL,
  T16_CS,
  T16_CB,
  T16_CJ
} t_format_16_sel;

// register width
typedef enum logic [3:0] {
  T16_W,
  T16_D,
  T16_Q
} t_format_16_wdh;

function logic signed [16:0] imm16 (t_format_16 i, t_format_16_sel sel, t_format_16_wdh wdh);
  logic [15:0] imm16 = '0;
  case (sel)
    T16_CR:
	imm16 = 'x;
    T16_CI:
      case (wdh)
        T16_W: {imm16[5], {imm16[4:2], imm16[7:6]}} = {i.ci.imm_12_12, i.ci.imm_06_02};
        T16_D: {imm16[5], {imm16[4:3], imm16[8:6]}} = {i.ci.imm_12_12, i.ci.imm_06_02};
        T16_Q: {imm16[5], {imm16[4:4], imm16[9:6]}} = {i.ci.imm_12_12, i.ci.imm_06_02};
	default: imm16 = 'x;
      endcase
    T16_CSS:
      case (wdh)
        T16_W: {imm16[5:2], imm16[7:6]} = i.css.imm_12_07;
        T16_D: {imm16[5:3], imm16[8:6]} = i.css.imm_12_07;
        T16_Q: {imm16[5:4], imm16[9:6]} = i.css.imm_12_07;
	default: imm16 = 'x;
      endcase
    T16_CIW:
      {imm16[5:4], imm[9:6], imm[2], imm[3]} = i.ciw.imm_16_05;
    T16_CL,
    T16_CS:
      case (wdh)
        T16_W: {imm16[5:3], imm16[2], imm16[  6]} = {i.cl.imm_12_10, i.cl.imm_06_05};
        T16_D: {imm16[5:3],           imm16[7:6]} = {i.cl.imm_12_10, i.cl.imm_06_05};
        T16_Q: {imm16[5:4], imm16[8], imm16[7:6]} = {i.cl.imm_12_10, i.cl.imm_06_05};
	default: imm16 = 'x;
      endcase
    T16_CJ:
      {imm16[11], imm16[4], imm16[9:8], imm16[10], imm16[6], imm16[7], imm16[3:1], imm16[5]} = i.cj.target;
    T16_CB:
      {imm16[8], imm16[4:3], imm16[7:6], imm16[2:1], imm16[5]} = {i.cb.off_12_10, i.cb.off_06_02};
    default: imm16 = 'x;
  endcase
endfunction: imm16

function logic [4:0] reg_5 (logic [2:0] reg_3);
  reg_5 = {2'b01, reg_3};
endfunction: reg_5

function ctli_t dec16 (frm16_t op, isa_t isa, int unsigned xw);
casez (op)
//  fedc_ba98_7654_3210                pc,     rs1,     rs2,                 imm,     alu,     br,   st,ste,    ld,lde,     wb,wbe,   csr,ill
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,                  'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b000?_????_????_??00: dec32 = '{PC_PC2, A1_SP , A2_IMM, 4*imm16(op,T16_CIW), AO_ADD,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, ~|imm16(op,T16_CIW)}; // C.ADDI4SP
16'b000?_????_????_??00: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction
16'b0000_0000_0000_0000: dec32 = '{PC_PC2,      'x,      'x,    'x,      'x,     'x,   'x, '0,    'x, '0,     'x, '0,    'x, '1}; // illegal instruction

32'b????_????_????_????_????_????_?001_0111: dec32 = '{PC_PC4, A1_PC , A2_IMM, IMM_U, AO_ADD,     'x,   'x, '0,    'x, '0, WB_ALU, '1, CSR_N, '0};  // auipc
32'b????_????_????_????_????_????_?110_1111: dec32 = '{PC_ALU, A1_PC , A2_IMM, IMM_J, AO_ADD,     'x,   'x, '0,    'x, '0, WB_PC4, '1, CSR_N, '0};  // jal
32'b????_????_????_????_?000_????_?110_0111: dec32 = '{PC_ALU, A1_RS1, A2_IMM, IMM_I, AO_ADD,     'x,   'x, '0,    'x, '0, WB_PC4, '1, CSR_N, '0};  // jalr
endcase
endfunction: dec16

endpackage: riscv_isa_pkg
