import riscv_isa_pkg::*;

module r5p_muldiv #(
  int unsigned XW = 32
)(
  // control
  input  ctl_m_t        ctl,
  // data input/output
  input  logic [XW-1:0] rs1,  // source register 1
  input  logic [XW-1:0] rs2,  // source register 2
  output logic [XW-1:0] rd    // destination register
);

// minux max (most negative value)
localparam logic [XW-1:0] M8 = {1'b1, {XW-1{1'b0}}};
// minus 1 (-1)
localparam logic [XW-1:0] M1 = '1;

logic [2-1:0][XW-1:0] mul;
logic        [XW-1:0] div;
logic        [XW-1:0] rem;

// NOTE:
// for signed*unsigned multiplication to work,
// the first operand must be sign extended to the LHS (result) width

// multiplication
always_comb
case (ctl.s12) inside
  2'b00  : mul = 64'($unsigned(rs1)) * $unsigned(rs2);
  2'b10  : mul = 64'(  $signed(rs1)) * $unsigned(rs2);
  2'b11  : mul = 64'(  $signed(rs1)) *   $signed(rs2);
  default: mul = 'x;
endcase

// division
always_comb
case (ctl.s12) inside
  2'b00  : div = ~|rs2 ? '1 :                            $unsigned(rs1) / $unsigned(rs2);
  2'b11  : div = ~|rs2 ? '1 : (rs1==M8 & rs2==M1) ? M8 :   $signed(rs1) /   $signed(rs2);
  default: div = 'x;
endcase

// reminder
always_comb
case (ctl.s12) inside
  2'b00  : rem = ~|rs2 ? rs1 :                            $unsigned(rs1) / $unsigned(rs2);
  2'b11  : rem = ~|rs2 ? rs1 : (rs1==M8 & rs2==M1) ? '0 :   $signed(rs1) /   $signed(rs2);
  default: rem = 'x;
endcase

always_comb
case (ctl.op) inside
  M_MUL: rd = mul[0];
  M_MUH: rd = mul[1];
  M_DIV: rd = div;
  M_REM: rd = rem;
endcase

logic unsigned [2*XW-1:0] mul64u;
logic   signed [2*XW-1:0] mul64s;

assign mul64u =   $signed(rs1) * $unsigned(rs2);
assign mul64s =   $signed(rs1) * $unsigned(rs2);

endmodule: r5p_muldiv