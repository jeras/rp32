../../../src/mem_if.vh